/*
 * simple なサンプル
 *
 * このサンプルは tecsgen/test/simple 階層に置いて実行する
 * Linux, Cygwin 環境で実行できるはず
 */

import_C( "tecs.h" );
import( <cygwin_kernel.cdl> );
import( <tSysLog.cdl> );

/* SysLog */
cell tSysLog SysLog {};

/* Kernel */
cell tKernel Kernel {};

/* typedef int32_t ER; */

namespace nMySpace {
	signature sSimple {
		ER  func1( [in]int32_t inval );
		ER  func2( [out,string]char_t *str );
	};

	celltype tSimpleServer {
		entry sSimple eEnt;
	};

	celltype tSimpleClient {
		call sSimple cCall;
	};
};

region rServer {
	cell nMySpace::tSimpleServer SimpleServer {
	};
};

[to_through(rServer)]
region rClient {
	cell nMySpace::tSimpleClient SimpleClient {
		[through(TLVTracePlugin,"")]
			cCall = rServer::SimpleServer.eEnt;
	};
};
