/*
 *  @(#) $Id: target_syssvc_inst.cdl 109 2008-05-28 14:33:39Z ertl-hiro $
 */

/*
 *		�������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ��Ⱦ夲����
 *		��Skyeye�ѡ�
 */

/*
 *  �ʰ�SIO�ɥ饤�Ф��Ȥ߾夲����
 */
cell tSerialPort SerialPort1;


cell tSIOPortSkyeye SIOPortTarget{
	ciSIOCBR = SerialPort1.eiSIOCBR;
};

/*
 *  �����ƥ�������٥���Ϥ��Ⱦ夲����
 */
cell tPutLogSkyeye PutLogTarget {
	cSIOPort = SIOPortTarget.eSIOPort;
};

