/*
 *  @(#) $Id: tLogTask.cdl 426 2009-07-17 05:06:29Z ertl-takuya $
 */

/*
 *		�����ƥ���������Υ���ݡ��ͥ�ȵ��ҥե�����
 */

signature sLogTask {
	ER		flush([in] uint_t count);
};

[singleton]
celltype tLogTaskMain{
	entry sTaskBody		eLogTaskBody;
	entry sLogTask		eLogTask;
	call sSerialPort	cSerialPort;	/* ���ꥢ��ɥ饤�ФȤ���³ */
	call snSerialPort	cnSerialPort;	/* ���ꥢ��ɥ饤�д����Ȥ���³ */
	call sSysLog		cSysLog;		/* �����ƥ����ǽ�Ȥ���³ */
	call sPutLog		cPutLog;		/* ���٥���ϤȤ���³ */

	attr {
		RELTIM	interval = 10;			/* ��������ư��ֳ� */
		RELTIM	flushWait = 1;			/* �ե�å����Ԥ���ñ�̻��� */
	};
	factory {
		write("tecsgen.cfg", "ATT_TER({ TA_NULL, 0, tLogTask_terminate });");
	};
	FACTORY {
		write("tecsgen.cfg", "#include \"syssvc/tLogTask.h\"");
	};
};
[singleton,active]
composite tLogTask{
	entry sTaskBody		eLogTaskBody;
	entry sTask       	eTask;	/* ���������ʥ���������ƥ������ѡ�*/
	entry siTask    	eiTask;	/* �����������󥿥�������ƥ������ѡ�*/
    [optional] call	sTaskExceptionBody	cExceptionBody;

	entry sLogTask		eLogTask;
	
	call sSerialPort	cSerialPort;	/* ���ꥢ��ɥ饤�ФȤ���³ */
	call snSerialPort	cnSerialPort;	/* ���ꥢ��ɥ饤�д����Ȥ���³ */
	call sSysLog		cSysLog;		/* �����ƥ����ǽ�Ȥ���³ */
	call sPutLog		cPutLog;		/* ���٥���ϤȤ���³ */

	attr {
		[omit] ATR		taskAttribute = C_EXP("TA_NULL");
		[omit] ATR		exceptionAttribute= C_EXP("TA_NULL");
		[omit] PRI  	priority;			/* �������ν��ͥ���� */
		[omit] SIZE 	stackSize;			/* �������Υ����å������� */
		RELTIM	interval = 10;			/* ��������ư��ֳ� */
		RELTIM	flushWait = 1;			/* �ե�å����Ԥ���ñ�̻��� */
	};
	cell tLogTaskMain LogTaskMain{
		/* �ƤӸ� */
		cSerialPort  => composite.cSerialPort;
		cnSerialPort => composite.cnSerialPort;
		cSysLog      => composite.cSysLog;
		cPutLog      => composite.cPutLog;
		/* °�� */
		interval     =  composite.interval;
		flushWait   =  composite.flushWait;
	};
	cell tTask Task{
		/* �ƤӸ� */
		cBody         =  LogTaskMain.eLogTaskBody;
		cExceptionBody=> composite.cExceptionBody;
		/* °�� */
		taskAttribute = composite.taskAttribute;
		exceptionAttribute = composite.exceptionAttribute;
		priority      = composite.priority;
		stackSize    = composite.stackSize;
	};
	/* ������ */
	composite.eLogTaskBody => LogTaskMain.eLogTaskBody;
	composite.eLogTask     => LogTaskMain.eLogTask;
	composite.eTask        => Task.eTask;
	composite.eiTask       => Task.eiTask;
};

