/*
 * 
 */
signature sPutLog {
	void	putChar([in] char c);
};

[singleton]
celltype tPutLogSkyeye {
	entry sPutLog	ePutLog;
	call  sSIOPort  cSIOPort;
};
