 /*
  * ���¸�����󶡤���ؿ�
  */
signature sSIOPort {
 	void	open(void);
	void	close(void);
	bool_t	putChar([in] char c);
	int_t	getChar(void);
	void	enableCBR([in] uint_t cbrtn);
	void	disableCBR([in] uint_t cbrtn);
};
/*
 * ���¸���ؤΥ�����Хå�
 */
signature siSIOCBR {
	void	readySend(void);
	void	readyReceive(void);
};

/* ������Хå��롼����μ����ֹ� */
const uint_t SIO_RDY_SND = 1;		/* ������ǽ������Хå� */
const uint_t SIO_RDY_RCV = 2;		/* �������Υ�����Хå� */

celltype tSIOPortSkyeyeMain {
	entry sSIOPort	eSIOPort;
	call siSIOCBR	ciSIOCBR;

	entry sInitializeRoutineBody eInitialize; /* ��������� */
	entry sTerminateRoutineBody eTerminate;   /* ��λ���� */

	entry siHandlerBody eiISR;/* ����ߥ����ӥ��롼���� */
	
	attr {
		/*Skyeye�ѤΥ��ɥ쥹*/
		uint32_t  uartBase;
	};
	var {
		/*
		 * skyeye��
		 */
		bool_t	openFlag;			/* �����ץ�Ѥߥե饰 */
		bool_t	receiveFlag;			/* ����ʸ���Хåե�ͭ���ե饰 */
		char	receiveBuffer;			/* ����ʸ���Хåե� */
		bool_t	receiveReady;			/* �������Υ�����Хå����ĥե饰 */
		/* SkyEye�ξ��������Ͼ�ˤǤ���Τǡ�����ʸ���Хåե���ɬ�פʤ� */
     	bool_t	sendReady;			/* �������Υ�����Хå����ĥե饰 */
	};
	FACTORY {
		write("$ct$_factory.h", "#include \"at91skyeye.h\"");
	};
};

[active]
composite tSIOPortSkyeye {
	entry sSIOPort	eSIOPort;
	call siSIOCBR	ciSIOCBR;

	attr {
		/*Skyeye�ѤΥ��ɥ쥹*/
		//uint32_t* uartBase = C_EXP("(USART0_BASE)");
		uint32_t uartBase = 0xFFFD0000;
	};

	cell tSIOPortSkyeyeMain SIOPortMain {
		ciSIOCBR => composite.ciSIOCBR;
		uartBase = composite.uartBase;
	};
	/*
	 *  �ʰ�SIO�ɥ饤�Фν���������롼����
	 */
	cell tInitializeRoutine InitializeSIO{
		cInitializeRoutine = SIOPortMain.eInitialize;
	};
	/*
	 *  �ʰ�SIO�ɥ饤�Фν�λ�����롼����
	 */
	cell tTerminateRoutine TerminateSIO{
		cTerminateRoutine = SIOPortMain.eTerminate;
	};
	cell tISRWithConfigInterrupt SIOPortSkyeyeISR{
		ciBody =  SIOPortMain.eiISR;
		interruptNumber   =  2;
		interruptPriority = -2;
	};
	composite.eSIOPort => SIOPortMain.eSIOPort;
};
	