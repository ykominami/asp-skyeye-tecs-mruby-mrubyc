/*
 *  @(#) $Id: target_syssvc_decl.cdl 109 2008-05-28 14:33:39Z ertl-hiro $
 */

/*
 *		�������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ������Skyeye�ѡ�
 */

/*
 *  �ʰ�SIO�ɥ饤�Ф����
 */
import("tSIOPortSkyeye.cdl");

/*
 *  �����ƥ�������٥���Ϥ����
 */
import("tPutLogSkyeye.cdl");

/*
 *  ���������Υ����å�������
 */
const uint_t LogTaskStackSize = 131072;
