/* 
/*
 * mruby Bridge  
 * $Id: Sample.cdl 1846 2012-11-11 02:35:54Z ritsumei-takuya $
 *
 * 
 *
 *  +----------------------------------+           +---------------------+          +-------------+
 *  | mruby object                     |           |                     |          |             |
 *  |taskBridge=                       |  sTask    |  tMrubyBridgesTask  |  sTask   |   tTask     |
 *  | TMrubyBridgesTask("TaskBridge")  |==========>|     TaskBridge      |----------|> MainTask   |
 *  |                                  |  �δؿ��� |                     |cCall eEnt|             |
 *  |                                  |           |                     |          |             |
 *  +----------------------------------+           +---------------------+          +-------------+
 *
 *�������˥��㵭��
 *
 *   sTask �� �ؿ����󥿥ե����������
 *            �����Ȥ�����Ƭʸ�� s ���ղä���
 * 
 *    �����˥��� sTask�ˤ�activate(��������ư)�ʤɥ�����������
 *
 *�����륿���׵���
 *
 *   tMrubyBridgesTask �� �֥�å�����Υ��륿���� (MrubyBridgePlugin �ˤ������)
 *   tTask             �� �Ƥ���Υ��륿����
 *
 */
/*
 *  �����ͥ륪�֥������Ȥ����
 */
import(<kernel.cdl>);

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ����
 */
import(<target_syssvc_decl.cdl>);

/*
 *  ���ꥢ��ɥ饤�Ф����
 */
import(<syssvc/tSerialPort.cdl>);

/*
 *  �����ƥ����ǽ�����
 */
import(<syssvc/tSysLog.cdl>);

/*
 *  �����ƥ�������������
 */
import(<syssvc/tLogTask.cdl>);

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ��Ȥ߾夲����
 */
import(<target_syssvc_inst.cdl>);

/* mruby������ */
import(<tMruby.cdl>);

/*
 *  �Ȥ߾夲����
 */

cell nMruby::tMruby Mruby{
	mrubyFile="mrb_sample_kernel_obj.rb";
	cSerialPort = SerialPort1.eSerialPort;
};


cell tSerialPort SerialPort1 {
	/* �ƤӸ��η�� */
	cSIOPort = SIOPortTarget.eSIOPort;
	receiveBufferSize = 256;
	sendBufferSize = 256;
};

cell tSysLog SysLog {
	/* �ƤӸ��η�� */
	cPutLog = PutLogTarget.ePutLog;
	logBufferSize = 32;
};

cell tLogTask LogTask {
	/* �ƤӸ��η�� */
	cSerialPort = SerialPort1.eSerialPort;
	cnSerialPort = SerialPort1.enSerialPort;
	cSysLog = SysLog.eSysLog;
	cPutLog = PutLogTarget.ePutLog;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = 3;
	stackSize = LogTaskStackSize;
	
};

cell tKernel ASPKernel{
};

cell tTask MrubyTask {
	/* �ƤӸ��η�� */
	cBody = Mruby.eMrubyBody;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = C_EXP("MAIN_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};

/*
 * �����˥���ץ饰���� MrubyBridgePlugin �θƤӽФ���
 *
 * MrubyBridgePlugin �ˤ��
 * ���֥�å��Υ��륿���� tMrubyBridgesTask ������� 
 *   gen/tmp_MrubyBridgePlugin_0.cdl ����������롣
 *   sTask ����ʬ�ϡ������˥���̾��
 * �����륿���ץ����� gen/nMruby_STask.c �ˡ�mruby �� 
 *   TMrubyBridgesTask ���饹��������ɤ���������롣
 */

/*
 * �֥�å����������
 *
 * mruby ���顢TMrubyBridgesTask ���饹�� Bridge �Ȥ��ƻ��Ȥ���롣
 *   ex) taskBridge = TECS::STask.new "TaskBridge"
 *
 * cTECS �� signature�����ʤ�� sTask �δؿ�����STask
 * �Υ��󥹥��󥹥᥽�åɤȤ���������졢�ƤӽФ����Ȥ��Ǥ��롣
 *   ex) taskBridge.activate
 */

celltype tTaskBody{
	entry sTaskBody eTaskBody;
};

cell tTaskBody MainTaskBody{
};

cell tTask MainTask {
	/* �ƤӸ��η�� */
	cBody = MainTaskBody.eTaskBody;
	/* °�������� */
	priority = 1;
	stackSize = C_EXP("STACK_SIZE");
};
//generate( MrubyBridgePlugin, sTask, "include=activate" );
generate( MrubyBridgePlugin, sTask, "" );
cell nMruby::STask TaskBridge {
	cTECS = MainTask.eTask;
};
