/*
 *		����ץ�ץ����(1)�Υ���ݡ��ͥ�ȵ��ҥե�����
 */

/*
 *  �����ͥ륪�֥������Ȥ����
 */
import(<kernel.cdl>);

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ����
 */
import(<target_syssvc_decl.cdl>);

/*
 *  ���ꥢ��ɥ饤�Ф����
 */
import(<syssvc/tSerialPort.cdl>);

/*
 *  �����ƥ����ǽ�����
 */
import(<syssvc/tSysLog.cdl>);

/*
 *  �����ƥ�������������
 */
import(<syssvc/tLogTask.cdl>);

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ��Ȥ߾夲����
 */
import(<target_syssvc_inst.cdl>);

/* mruby������ */
import(<tMruby.cdl>);

/*
 * �����˥���ץ饰���� MrubyBridgePlugin �θƤӽФ���
 */
generate( MrubyBridgePlugin, sKernel, "" );



/*
 *  ����ץ�ץ��������
 */
	cell nMruby::tsKernel BridgeKernel {
		cTECS = ASPKernel.eKernel;
	};

	//Kernel
	cell tKernel ASPKernel{
	};

[singleton]
celltype tSample1 {
	require tKernel.eKernel;// �ƤӸ�̾�ʤ����㡧delay��
	//require cKernel = tKernel.eKernel;// �ƤӸ�̾������㡧cKernel_delay��
	require ciKernel = tKernel.eiKernel;// �ƤӸ�̾������㡧ciKernel_��

	call sTask          cTask;
    /*call sMrubyBody     cMrubyBody;*/

	call sSerialPort	cSerialPort;	/* ���ꥢ��ɥ饤�ФȤ���³ */
	call sSysLog		cSysLog;		/* �����ƥ����ǽ�Ȥ���³ */
	
	entry sTaskBody		eMainTask;	  /* Main������ */
	entry sTaskExceptionBody	eSampleException;/* �������㳰�����롼���� */
};

/*
 *  �Ȥ߾夲����
 */

cell tSerialPort SerialPort1 {
	/* �ƤӸ��η�� */
	cSIOPort = SIOPortTarget.eSIOPort;
	receiveBufferSize = 256;
	sendBufferSize = 256;
};

cell tSysLog SysLog {
	/* �ƤӸ��η�� */
	cPutLog = PutLogTarget.ePutLog;
	logBufferSize = 32;
};

cell tLogTask LogTask {
	/* �ƤӸ��η�� */
	cSerialPort = SerialPort1.eSerialPort;
	cnSerialPort = SerialPort1.enSerialPort;
	cSysLog = SysLog.eSysLog;
	cPutLog = PutLogTarget.ePutLog;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = 3;
	stackSize = LogTaskStackSize;
	
};

cell tTask MainTask {
	/* �ƤӸ��η�� */
	cBody = Sample1.eMainTask;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = C_EXP("MAIN_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};

cell tSample1 Sample1 {
	/* �ƤӸ��η�� */
	cTask =MainTask.eTask;

	cSerialPort = SerialPort1.eSerialPort;
	cSysLog = SysLog.eSysLog;
};

cell tTask MrubyTask0 {
	/* �ƤӸ��η�� */
	cBody = Mruby0.eMrubyBody;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = C_EXP("MID_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};

cell tTask MrubyTask2 {
	/* �ƤӸ��η�� */
	cBody = Mruby2.eMrubyBody;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = C_EXP("LOW_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};

cell nMruby::tMruby Mruby2{
	mrubyFile="mrb2.rb mrb21.rb";
	/* cSerialPort = SerialPort1.eSerialPort;*/
	cInit = VM_TECSInitializer.eInitialize;
    ida = 2;
};

cell nMruby::tMruby Mruby0{
	mrubyFile="mrb0.rb";
	/* cSerialPort = SerialPort1.eSerialPort;*/
	cInit = VM_TECSInitializer.eInitialize;
    ida = 0;
};


