/*
 *  @(#) $Id: tSerialPort.cdl 439 2009-07-22 09:08:30Z ertl-takuya $
 */

/*
 *		���ꥢ�륤�󥿥ե������ɥ饤�ФΥ���ݡ��ͥ�ȵ��ҥե�����
 */

typedef struct {
	uint_t		reacnt;				/* �����Хåե����ʸ���� */
	uint_t		wricnt;				/* �����Хåե����ʸ���� */
} T_SERIAL_RPOR;

signature sSerialPort {
	ER		open(void);
	ER		close(void);
	ER_UINT	read([out,size_is(length)] char *buffer, [in] uint_t length);
	ER_UINT	write([in,size_is(length)] const char *buffer, [in] uint_t length);
	ER		control([in] uint_t ioControl);
	ER		refer([out] T_SERIAL_RPOR *pk_rpor);
};

signature snSerialPort {
	bool_t	getChar([out] char *p_char);
};

/* ���ꥢ�륤�󥿥ե������ɥ饤�Ф�ư�������ѤΤ������� */
const uint_t IOCTL_NULL	= 0;		/* ����ʤ� */
const uint_t IOCTL_ECHO	= 0x0001;	/* ��������ʸ���򥨥����Хå� */
const uint_t IOCTL_CRLF	= 0x0010;	/* LF��������������CR���ղ� */
const uint_t IOCTL_FCSND = 0x0100;	/* �������Ф��ƥե������Ԥ� */
const uint_t IOCTL_FCANY = 0x0200;	/* �ɤΤ褦��ʸ���Ǥ������Ƴ� */
const uint_t IOCTL_FCRCV = 0x0400;	/* �������Ф��ƥե������Ԥ� */

celltype tSerialPortMain {
	entry sSerialPort	eSerialPort;
	entry snSerialPort	enSerialPort;

 	call sSIOPort		cSIOPort;	/* �ʰ�SIO�ɥ饤�ФȤ���³ */
	entry siSIOCBR		eiSIOCBR;
	
	call sSemaphore  cSendSemaphore;
	call siSemaphore ciSendSemaphore;

	call sSemaphore  cReceiveSemaphore;
	call siSemaphore ciReceiveSemaphore;
	
	attr {
		uint_t	receiveBufferSize = 256;	/* �����Хåե������� */
		uint_t	sendBufferSize = 256;	/* �����Хåե������� */
	};
	var {
		bool_t	openFlag = C_EXP("false");	/* �����ץ�Ѥߥե饰 */
		bool_t	errorFlag;			/* ���顼�ե饰 */
		uint_t	ioControl;				/* ư������������� */

		[size_is(receiveBufferSize)] char	*receiveBuffer;	/* �����Хåե� */
		uint_t	receiveReadPointer;		/* �����Хåե��ɽФ��ݥ��� */
		uint_t	receiveWritePointer;		/* �����Хåե�����ߥݥ��� */
		uint_t	receiveCount;			/* �����Хåե����ʸ���� */
		char	receiveFlowControl;			/* ����٤�START/STOP */
		bool_t	receiveStopped;		/* STOP�����ä����֤��� */

		[size_is(sendBufferSize)] char	*sendBuffer;	/* �����Хåե� */
		uint_t	sendReadPointer;		/* �����Хåե��ɽФ��ݥ��� */
		uint_t	sendWritePointer;		/* �����Хåե�����ߥݥ��� */
		uint_t	sendCount;			/* �����Хåե����ʸ���� */
		bool_t	sendStopped;		/* STOP�������ä����֤��� */
	};
};

composite tSerialPort{
	entry sSerialPort	eSerialPort;
	entry snSerialPort	enSerialPort;

 	call sSIOPort		cSIOPort;	/* �ʰ�SIO�ɥ饤�ФȤ���³ */
	entry siSIOCBR		eiSIOCBR;
	
	attr {
		uint_t	receiveBufferSize = 256;	/* �����Хåե������� */
		uint_t	sendBufferSize = 256;	/* �����Хåե������� */
	};
	/* �����ѤΥ��ޥե� */
	cell tSemaphore ReceiveSemaphore{
		attribute = C_EXP("TA_NULL");
		count = 0;
		max =1;
	};
	/* �����ѤΥ��ޥե� */
	cell tSemaphore SendSemaphore{
		attribute = C_EXP("TA_NULL");
		count = 1;
		max =1;
	};
	/* ���ꥢ��ݡ��Ȥ������� */
	cell tSerialPortMain SerialPortMain{
		/* �ƤӸ��η�� */
		cReceiveSemaphore  = ReceiveSemaphore.eSemaphore;
		ciReceiveSemaphore = ReceiveSemaphore.eiSemaphore;
		cSendSemaphore  = SendSemaphore.eSemaphore;
		ciSendSemaphore = SendSemaphore.eiSemaphore;
		/* �ƤӸ��Υ������ݡ��� */
		cSIOPort => composite.cSIOPort;
		/* °�� */
		receiveBufferSize = composite.receiveBufferSize;
		sendBufferSize = composite.sendBufferSize;
	};
	/* ������ */
	composite.eSerialPort  => SerialPortMain.eSerialPort;
	composite.enSerialPort => SerialPortMain.enSerialPort;
	composite.eiSIOCBR     => SerialPortMain.eiSIOCBR;
};
