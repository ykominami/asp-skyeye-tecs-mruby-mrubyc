/*
 *		����ץ�ץ����(1)�Υ���ݡ��ͥ�ȵ��ҥե�����
 */

/*
 *  �����ͥ륪�֥������Ȥ����
 */
import(<kernel.cdl>);

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ����
 */
import(<target_syssvc_decl.cdl>);

/*
 *  ���ꥢ��ɥ饤�Ф����
 */
import(<syssvc/tSerialPort.cdl>);

/*
 *  �����ƥ����ǽ�����
 */
import(<syssvc/tSysLog.cdl>);

/*
 *  �����ƥ�������������
 */
import(<syssvc/tLogTask.cdl>);

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ��Ȥ߾夲����
 */
import(<target_syssvc_inst.cdl>);

/* mruby������ */
import(<tMruby.cdl>);

/*
 *  ����ץ�ץ��������
 */
/*[singleton]
celltype tSample {
	require tKernel.eKernel;// �ƤӸ�̾�ʤ����㡧delay��
	//require cKernel = tKernel.eKernel;// �ƤӸ�̾������㡧cKernel_delay��
	require ciKernel = tKernel.eiKernel;// �ƤӸ�̾������㡧ciKernel_��
	call sTask          cTask;
    call sMrubyBody     cMrubyBody;

  
	call sSerialPort	cSerialPort;	// ���ꥢ��ɥ饤�ФȤ���³ 
	call sSysLog		cSysLog;		// �����ƥ����ǽ�Ȥ���³ 
	
	entry sTaskBody		eMainTask;	  // Main������ 
};
*/
/*
 *  �Ȥ߾夲����
 */


cell nMruby::tMruby Mruby{
	mrubyFile="mrb_sample.rb";
	cSerialPort = SerialPort1.eSerialPort;
};


cell tSerialPort SerialPort1 {
	/* �ƤӸ��η�� */
	cSIOPort = SIOPortTarget.eSIOPort;
	receiveBufferSize = 256;
	sendBufferSize = 256;
};

cell tSysLog SysLog {
	/* �ƤӸ��η�� */
	cPutLog = PutLogTarget.ePutLog;
	logBufferSize = 32;
};

cell tLogTask LogTask {
	/* �ƤӸ��η�� */
	cSerialPort = SerialPort1.eSerialPort;
	cnSerialPort = SerialPort1.enSerialPort;
	cSysLog = SysLog.eSysLog;
	cPutLog = PutLogTarget.ePutLog;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = 3;
	stackSize = LogTaskStackSize;
	
};

cell tKernel ASPKernel{
};

cell tTask MrubyTask1 {
	/* �ƤӸ��η�� */
	cBody = Mruby.eMrubyBody;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = C_EXP("MAIN_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};


cell tTask MrubyTask2 {
	/* �ƤӸ��η�� */
	cBody = Mruby2.eMrubyBody;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = C_EXP("MAIN_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};


cell nMruby::tMruby Mruby2{
	mrubyFile= "mrb_sample2.rb";
	cSerialPort = SerialPort1.eSerialPort;
};