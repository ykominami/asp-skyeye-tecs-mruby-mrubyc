/*
 *  @(#) $Id: tSysLog.cdl 1146 2010-10-13 07:36:12Z ritsumei-takuya $
 */

/*
 *		�����ƥ����ǽ�Υ���ݡ��ͥ�ȵ��ҥե�����
 */
import_C("t_syslog.h");

signature sSysLog {
	ER		write([in] uint_t priority, [in] const SYSLOG *p_syslog);
	ER_UINT	read([out] SYSLOG *p_syslog);
	ER		mask([in] uint_t logMask, [in] uint_t lowMask);
	ER		refer([out] T_SYSLOG_RLOG *pk_rlog);
};

[singleton]
celltype tSysLog {
	entry sSysLog	eSysLog;
	call sPutLog	cPutLog;		/* ���٥���ϤȤ���³ */

	attr {
		uint_t	logBufferSize;			/* ���Хåե������� */
	};
	var {
		[size_is(logBufferSize)] SYSLOG	*logBuffer;	/* ���Хåե� */
		uint_t	count = 0;			/* ���Хåե���Υ��ο� */
		uint_t	head = 0;			/* ��Ƭ�Υ��γ�Ǽ���� */
		uint_t	tail = 0;			/* ���Υ��γ�Ǽ���� */
		uint_t	lost = 0;			/* ����줿���ο� */
		uint_t	logMask = 0;		/* ���Хåե��˵�Ͽ���٤������� */
		uint_t	lowMaskNot = 0;     /* ���٥���Ϥ��٤������� */
	};
	FACTORY {
		/*
         * Syslog�����Ѥ������Makefile�����
		 */
		write("Makefile.tecsgen", "USE_SYSLOG = ture");
	};
};
