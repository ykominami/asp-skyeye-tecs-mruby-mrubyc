/*
 *		����ץ�ץ����(1)�Υ���ݡ��ͥ�ȵ��ҥե�����
 */

/*
 *  �����ͥ륪�֥������Ȥ����
 */
import(<kernel.cdl>);

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ����
 */
import(<target_syssvc_decl.cdl>);

/*
 *  ���ꥢ��ɥ饤�Ф����
 */
import(<syssvc/tSerialPort.cdl>);

/*
 *  �����ƥ����ǽ�����
 */
import(<syssvc/tSysLog.cdl>);

/*
 *  �����ƥ�������������
 */
import(<syssvc/tLogTask.cdl>);

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ��Ȥ߾夲����
 */
import(<target_syssvc_inst.cdl>);

/* mruby������ */
import(<tMruby.cdl>);

/*
 *  ����ץ�ץ��������
 */
[singleton]
celltype tSample1 {
	require tKernel.eKernel;// �ƤӸ�̾�ʤ����㡧delay��
	//require cKernel = tKernel.eKernel;// �ƤӸ�̾������㡧cKernel_delay��
	require ciKernel = tKernel.eiKernel;// �ƤӸ�̾������㡧ciKernel_��

	call sTask          cTask;
    /*call sMrubyBody     cMrubyBody;*/

	call sSerialPort	cSerialPort;	/* ���ꥢ��ɥ饤�ФȤ���³ */
	call sSysLog		cSysLog;		/* �����ƥ����ǽ�Ȥ���³ */
	
	entry sTaskBody		eMainTask;	  /* Main������ */
	entry sTaskExceptionBody	eSampleException;/* �������㳰�����롼���� */
};

/*
 *  �Ȥ߾夲����
 */

cell tSerialPort SerialPort1 {
	/* �ƤӸ��η�� */
	cSIOPort = SIOPortTarget.eSIOPort;
	receiveBufferSize = 256;
	sendBufferSize = 256;
};

cell tSysLog SysLog {
	/* �ƤӸ��η�� */
	cPutLog = PutLogTarget.ePutLog;
	logBufferSize = 32;
};

cell tLogTask LogTask {
	/* �ƤӸ��η�� */
	cSerialPort = SerialPort1.eSerialPort;
	cnSerialPort = SerialPort1.enSerialPort;
	cSysLog = SysLog.eSysLog;
	cPutLog = PutLogTarget.ePutLog;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = 3;
	stackSize = LogTaskStackSize;
	
};

cell tKernel ASPKernel{
};

cell tTask MainTask {
	/* �ƤӸ��η�� */
	cBody = Sample1.eMainTask;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = C_EXP("MAIN_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};

cell tSample1 Sample1 {
	/* �ƤӸ��η�� */
	cTask =MainTask.eTask;

	cSerialPort = SerialPort1.eSerialPort;
	cSysLog = SysLog.eSysLog;
};
