/*
 *		����ץ�ץ����(1)�Υ���ݡ��ͥ�ȵ��ҥե�����
 */

/*
 *  �����ͥ륪�֥������Ȥ����
 */
import("kernel.cdl");

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ����
 */
import("target_syssvc_decl.cdl");

/*
 *  ���ꥢ��ɥ饤�Ф����
 */
import("syssvc/tSerialPort.cdl");

/*
 *  �����ƥ����ǽ�����
 */
import("syssvc/tSysLog.cdl");

/*
 *  �����ƥ�������������
 */
import("syssvc/tLogTask.cdl");

/*
 *  �������åȰ�¸�Υ����ƥॵ���ӥ�����ݡ��ͥ�Ȥ��Ȥ߾夲����
 */
import("target_syssvc_inst.cdl");

/*
 *  ����ץ�ץ��������
 */
[singleton]
celltype tSample1 {
	require tKernel.eKernel;// �ƤӸ�̾�ʤ����㡧delay��
	//require cKernel = tKernel.eKernel;// �ƤӸ�̾������㡧cKernel_delay��
	require ciKernel = tKernel.eiKernel;// �ƤӸ�̾������㡧ciKernel_��

	call sTask		    cTask[4];	/* ��������� */
	call sCyclic        cCyclic;
	call sAlarm         cAlarm;

	call sSerialPort	cSerialPort;	/* ���ꥢ��ɥ饤�ФȤ���³ */
	call sSysLog		cSysLog;		/* �����ƥ����ǽ�Ȥ���³ */
	
	entry sTaskBody		eMainTask;	  /* Main������ */
	entry sTaskBody		eSampleTask[3];/* �¹Լ¹Ԥ���륿���� */
	entry sTaskExceptionBody	eSampleException[3];/* �������㳰�����롼���� */
	
	entry siHandlerBody eiCyclicHandler;/* �����ϥ�ɥ�*/
	entry siHandlerBody eiAlarmHandler; /* ���顼��ϥ�ɥ� */
};

/*
 *  �Ȥ߾夲����
 */

cell tSerialPort SerialPort1 {
	/* �ƤӸ��η�� */
	cSIOPort = SIOPortTarget.eSIOPort;
	receiveBufferSize = 256;
	sendBufferSize = 256;
};

cell tSysLog SysLog {
	/* �ƤӸ��η�� */
	cPutLog = PutLogTarget.ePutLog;
	logBufferSize = 32;
};

cell tLogTask LogTask {
	/* �ƤӸ��η�� */
	cSerialPort = SerialPort1.eSerialPort;
	cnSerialPort = SerialPort1.enSerialPort;
	cSysLog = SysLog.eSysLog;
	cPutLog = PutLogTarget.ePutLog;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = 3;
	stackSize = LogTaskStackSize;
	
};

/* Sample1�Υץ�ȥ�������� */
cell tSample1 Sample1;


cell tKernel ASPKernel{
};

cell tTask MainTask {
	/* �ƤӸ��η�� */
	cBody = Sample1.eMainTask;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = C_EXP("MAIN_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};

cell tTask Task1 {
	/* �ƤӸ��η�� */
	cBody = Sample1.eSampleTask[0];
	cExceptionBody = Sample1.eSampleException[0];
	  /* °�������� */
	priority = C_EXP("MID_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};

cell tTask Task2 {
	/* �ƤӸ��η�� */
	cBody = Sample1.eSampleTask[1];
	cExceptionBody = Sample1.eSampleException[1];
	/* °�������� */
	priority = C_EXP("MID_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};

cell tTask Task3 {
	/* �ƤӸ��η�� */
	cBody = Sample1.eSampleTask[2];
	cExceptionBody = Sample1.eSampleException[2];
	/* °�������� */
	priority = C_EXP("MID_PRIORITY");
	stackSize = C_EXP("STACK_SIZE");
};

cell tCyclicHandler CyclicHandler {
	/* �ƤӸ��η�� */
	ciBody = Sample1.eiCyclicHandler;
	/* °�������� */
	cyclicTime = 2000;
};

cell tAlarmHandler AlarmHandler {
	ciBody = Sample1.eiAlarmHandler;
};

cell tSample1 Sample1 {
	/* �ƤӸ��η�� */
	cTask[ 0 ] =MainTask.eTask;
	cTask[ 1 ] =Task1.eTask;
	cTask[ 2 ] =Task2.eTask;
	cTask[ 3 ] =Task3.eTask;

	cCyclic = CyclicHandler.eCyclic;
	cAlarm  = AlarmHandler.eAlarm;

	cSerialPort = SerialPort1.eSerialPort;
	cSysLog = SysLog.eSysLog;
};
